../xschem/user_analog_project_wrapper.spice